module ALU (
    
);
    
endmodule