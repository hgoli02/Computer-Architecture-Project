module ALU_CONTROLLER(alu_operation, opcode, func, clk);

    output [3:0] alu_operation;
    reg [3:0] alu_operation;
    input [5:0] opcode;
    input [5:0] func;
    input clk;


    // R instructions
    if (opcode == 6'b000000) begin
        if(func == 6'b000000 || func == 6'b000100) //SLL, SLLV
            alu_operation = 4'd5;

        if(func == 6'b000010 || func == 6'b000110) //SRL, SRLV
            alu_operation = 4'd6;

        if(func == 6'b100110) //xor
            alu_operation = 4'd1;

        if(func == 6'b100010) // sub
            alu_operation = 4'd10;

        if(func == 6'b101010) // slt
            alu_operation = 4'd7;

        if(func == 6'b100011) //sub unsigned
            alu_operation = 4'd11;

        if(func == 6'b100101) // OR
            alu_operation = 4'd2;

        if(func == 6'b100111) //NOR
            alu_operation = 4'd4;

        if(func == 6'b100001) //add unsigned
            alu_operation = 4'd8;

        if(func == 6'b011000) //mult
            alu_operation = 4'd12;

        if(func == 6'b011010) //div
            alu_operation = 4'd13;

        if(func == 6'b100100) //AND
            alu_operation = 4'd3;

        if(func == 6'b100000) //add
            alu_operation = 4'd9;

        
    end
    
    // I instructions
    else begin
        if(opcode == 6'b001110) //XORi
            alu_operation = 4'd1;

        if(opcode == 6'b001010) //SLTi
            alu_operation = 4'd7;

        if(opcode == 6'b001000) //ADDi
            alu_operation = 4'd8;

        if(opcode == 6'b001100) //ANDi
            alu_operation = 4'd3;

        if(opcode == 6'b001101) //ORi 
            alu_operation = 4'd2;   

         if(opcode == 6'b001001) //ADDiu (unsigned) 
            alu_operation = 4'd8;   
        end
endmodule
