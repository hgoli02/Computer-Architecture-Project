module LeftShifter #(parameter count = 1) (in, out);
    input 


endmodule