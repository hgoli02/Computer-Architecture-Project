module CU (
    ports
);
    
endmodule