module cache_controller (
    
);
    
endmodule