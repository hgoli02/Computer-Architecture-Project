module alu (
    
);
    
endmodule