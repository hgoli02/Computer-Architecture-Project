module cache (
    
);
    
endmodule